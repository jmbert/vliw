
`define SINGLE 	6'b000000
`define NOP	26'b0

`define LUI 	6'b000001

`define OPI_ART 6'b000010
`define ADDUI	4'b0000
`define XORUI	4'b0001
`define ANDUI	4'b0010
`define ORUI	4'b0011
