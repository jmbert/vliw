
`define SINGLE 	6'b000000
`define NOP	26'b0

`define LUI 	6'b000001
`define LUUI	1'b0
`define LSUI	1'b1

`define OPI_ART 6'b000010
`define ADDUI	4'b0000
`define XORUI	4'b0001
`define ANDUI	4'b0010
`define ORUI	4'b0011

`define JALR	6'b000100
`define JALRFN	3'b000

`define JAL	6'b000101
