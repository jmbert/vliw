
`define SINGLE 	6'b000000
`define NOP	26'b0

`define OPI_16 	6'b000001

`define LUUI	5'b00000
`define LSUI	5'b00001
